package tp1_pkg is

	type t_semaforo_state is (S0, S1, S2, S3, S4, S5);

end package;